******************** STL ver 2.3 T element basic model ********************

*** Notice *** ------------------------------------------------------*
* TエレメントによるSTL基本形（バス配線で寄生容量接続有り）のテンプレート

*--------------------------------------------------------------------*


*** STL Circuit *** -------------------------------------------------*

Vs1             101     0       PULSE( 0 2 1n 200p 200p 1.8n 4n )
Rin1            101     102     50

T1_STL_3        102     0       optpt1  0       Z0=50   TD=630.8p       $ LEN=100m
C1              optpt1  0       10p
T2_STL_8        optpt1  0       optpt2  0       Z0=50   TD=630.8p       $ LEN=100m
C2              optpt2  0       10p
T3_STL_3        optpt2  0       optpt3  0       Z0=50   TD=630.8p       $ LEN=100m

RT1             optpt3  0       50

*--------------------------------------------------------------------*


*** Versus Circuit *** ----------------------------------------------*

Vsvs1          1001    0       PULSE( 0 2 1n 200p 200p 1.8n 4n )
Rinvs1         1001    1002    50
Tvs1           1002    0       vspt1   0       z0=50   TD=630.8p
Tvs2           vspt1   0       vspt2   0       z0=50   TD=630.8p
Tvs3           vspt2   0       vspt3   0       z0=50   TD=630.8p
RTvs1          vspt3   0       50

*--------------------------------------------------------------------*


*** Netlist Commands *** --------------------------------------------*

.WIDTH OUT=132
.TRAN 50p 40n 20n
.PRINT v(optpt1) v(optpt2) v(optpt3) v(vspt1) v(vspt2) v(vspt3)
.END

*--------------------------------------------------------------------*
